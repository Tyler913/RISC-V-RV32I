module ALU (
    input wire pll_1_200MHz,
    input wire pll_1_locked
);


endmodule
